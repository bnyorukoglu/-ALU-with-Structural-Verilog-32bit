module and_4input(S, A, B, C, D);

input   A,B,C, D;
output  S;

and and0(S, A, B, C, D);
endmodule